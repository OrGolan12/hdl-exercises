module comparator_1bit (
    input a,
    input b,
    output y
);

assign y = a & ~b;

endmodule

